//TODO - do all connections for TH here


