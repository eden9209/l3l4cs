`ifndef L3L4CS_DEFINES_SV
    `define L3L4CS_DEFINES_SV

    `define L3L4CS_TB       l3l4cs_tb
    `define L3L4CS_TH      `L3L4CS_TB.l3l4cs_th
    `define L3L4CS_TOP     `L3L4CS_TB.l3l4cs_top

    `define CS_AGENT_PER_L3L4CS_NUM 1
	`define AXI_AGENT_PER_L3L4CS_NUM 1
    `define AXI_WRPS_NUM 2

// ---------------------------------------------------------------------------
`endif // L3L4CS_DEFINES_SV

