   `include "uvm_macros.svh"

   import uvm_pkg::*;
   import gk_base_types_pkg::*;
   import gk_base_pkg::*;
   import ce_base_pkg::*;
   import ce_base_types_pkg::*;
   import gk_base_global_pkg::*;

   import axis_vwrp_pkg::*;
   import l3l4cs_global_pkg::*;

   import l3l4cs_axis_wrap_types_pkg::*;

   import l3l4cs_axis_wrap_pkg::*;
   import eth_p_agent_pkg::*;
   import eth_vip_pkg::*;


   import l3l4cs_cs_agent_pkg::*;
  

   import eth_vip_types_pkg::*;

   import l3l4cs_pkg::*;
   

  //  `include "direct/l3l4cs_frames_no_vlan_ipv4_tcp_test.sv"  
  //  `include "direct/l3l4cs_frames_no_vlan_ipv4_udp_test.sv"  
  //  `include "direct/l3l4cs_frames_with_vlan_ipv4_tcp_test.sv"  
  //  `include "direct/l3l4cs_frames_with_vlan_ipv4_udp_test.sv"  
  //  `include "direct/l3l4cs_length_error_test.sv"  
  //  `include "direct/l3l4cs_non_ip_test.sv"  
  //  `include "direct/l3l4cs_non_tcp_udp_test.sv"  

  //  `include "direct/l3l4cs_min_total_len_test.sv"  
  //  `include "direct/l3l4cs_max_total_len_jambo_test.sv"  

  //  `include "direct/l3l4cs_no_packet_recived_test.sv"  


    `include "random/l3l4cs_random_testing.sv"  
  // `include "direct/l3l4cs_corner_testing.sv"  
   `include "direct/l3l4cs_direct_testing.sv"  


 

