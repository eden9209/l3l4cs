`define CS_AGENT_DATA_WD 2
`define CS_AGENT_VLD_WD  1
// `define CS_AGENT_LANES 8
// `define CS_AGENT_DATA_WORD 10
 `define CS_AGENT_STREMAS 1

